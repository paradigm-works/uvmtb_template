//----------------------------------------------------------------------
// This File: CYCLE.sv
// Author:    cliff.cummings@paradigm-works.com
// SPDX-License-Identifier: MIT
//----------------------------------------------------------------------

`ifndef CYCLE
  `define CYCLE 10
`endif
`timescale 1ns/1ns
